library IEEE;
use IEEE.std_logic_1164.all;

entity ULA is

    port(

    );
    
    end ULA;

architecture comportamento of ULA is 

    begin
        --Fazer a ULA
    
    end comportamento;