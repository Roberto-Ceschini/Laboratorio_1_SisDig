--vou fazer o cdigo da and