library IEEE;
use IEEE.std_logic_1164.all;

entity complemento_2 is 

    port (

        num: in std_logic_vector (3 downto 0); --Entradas: numero a ser complementado
        saida: out std_logic_vector (3 downto 0) -- Saidas: numero complementado
    );

end complemento_2;

architecture comportamento of complemento_2 is -- Funcao: realiza o complemento a 2 de um numero

    begin
     --falta fazer a architeture
    end comportamento;